module Multiply16logic
(
input [15:0] A, B,
output [15:0][15:0] R
);

// assign R[15] = (A[15] & B[0]) + (A[14] & B[1]) + (A[13] & B[2]) + (A[12] & B[3]) + (A[11] & B[4]) + (A[10] & B[5]) + (A[9] & B[6]) + (A[8] & B[7]) + (A[7] & B[8]) + (A[6] & B[9]) + (A[5] & B[10]) + (A[4] & B[11]) + (A[3] & B[12]) + (A[2] & B[13]) + (A[1] & B[14]) + (A[0] & B[15]); 
// assign R[14] = (A[14] & B[0]) + (A[13] & B[1]) + (A[12] & B[2]) + (A[11] & B[3]) + (A[10] & B[4]) + (A[9] & B[5]) + (A[8] & B[6]) + (A[7] & B[7]) + (A[6] & B[8]) + (A[5] & B[9]) + (A[4] & B[10]) + (A[3] & B[11]) + (A[2] & B[12]) + (A[1] & B[13]) + (A[0] & B[14]);
// assign R[13] = (A[13] & B[0]) + (A[12] & B[1]) + (A[11] & B[2]) + (A[10] & B[3]) + (A[9] & B[4]) + (A[8] & B[5]) + (A[7] & B[6]) + (A[6] & B[7]) + (A[5] & B[8]) + (A[4] & B[9]) + (A[3] & B[10]) + (A[2] & B[11]) + (A[1] & B[12]) + (A[0] & B[13]);
// assign R[12] = (A[12] & B[0]) + (A[11] & B[1]) + (A[10] & B[2]) + (A[9] & B[3]) + (A[8] & B[4]) + (A[7] & B[5]) + (A[6] & B[6]) + (A[5] & B[7]) + (A[4] & B[8]) + (A[3] & B[9]) + (A[2] & B[10]) + (A[1] & B[11]) + (A[0] & B[12]);
// assign R[11] = (A[11] & B[0]) + (A[10] & B[1]) + (A[9] & B[2]) + (A[8] & B[3]) + (A[7] & B[4]) + (A[6] & B[5]) + (A[5] & B[6]) + (A[4] & B[7]) + (A[3] & B[8]) + (A[2] & B[9]) + (A[1] & B[10]) + (A[0] & B[11]);
// assign R[10] = (A[10] & B[0]) + (A[9] & B[1]) + (A[8] & B[2]) + (A[7] & B[3]) + (A[6] & B[4]) + (A[5] & B[5]) + (A[4] & B[6]) + (A[3] & B[7]) + (A[2] & B[8]) + (A[1] & B[9]) + (A[0] & B[10]); 
// assign R[9] = (A[9] & B[0]) + (A[8] & B[1]) + (A[7] & B[2]) + (A[6] & B[3]) + (A[5] & B[4]) + (A[4] & B[5]) + (A[3] & B[6]) + (A[2] & B[7]) + (A[1] & B[8]) + (A[0] & B[9]); 
// assign R[8] = (A[8] & B[0]) + (A[7] & B[1]) + (A[6] & B[2]) + (A[5] & B[3]) + (A[4] & B[4]) + (A[3] & B[5]) + (A[2] & B[6]) + (A[1] & B[7]) + (A[0] & B[8]);
// assign R[7] = (A[7] & B[0]) + (A[6] & B[1]) + (A[5] & B[2]) + (A[4] & B[3]) + (A[3] & B[4]) + (A[2] & B[5]) + (A[1] & B[6]) + (A[0] & B[7]);
// assign R[6] = (A[6] & B[0]) + (A[5] & B[1]) + (A[4] & B[2]) + (A[3] & B[3]) + (A[2] & B[4]) + (A[1] & B[5]) + (A[0] & B[6]);
// assign R[5] = (A[5] & B[0]) + (A[4] & B[1]) + (A[3] & B[2]) + (A[2] & B[3]) + (A[1] & B[4]) + (A[0] & B[5]);
// assign R[4] = (A[4] & B[0]) + (A[3] & B[1]) + (A[2] & B[2]) + (A[1] & B[3]) + (A[0] & B[4]);
// assign R[3] = (A[3] & B[0]) + (A[2] & B[1]) + (A[1] & B[2]) + (A[0] & B[3]);
// assign R[2] = (A[2] & B[0]) + (A[1] & B[1]) + (A[0] & B[2]);
// assign R[1] = (A[1] & B[0]) + (A[0] & B[1]);
// assign R[0] = (A[0] & B[0]);

assign R[0][15:0] = { (B[0] & A[15]) , (B[0] & A[14]) , (B[0] & A[13]) , (B[0] & A[12]) , (B[0] & A[11]) , (B[0] & A[10]) , (B[0] & A[9]) ,  (B[0] & A[8]) ,  (B[0] & A[7]) ,  (B[0] & A[6]) ,  (B[0] & A[5]) ,  (B[0] & A[4]) ,  (B[0] & A[3]) ,  (B[0] & A[2]) ,  (B[0] & A[1]) ,  (B[0] & A[0]) }; 
assign R[1][15:0] = { (B[1] & A[14]) , (B[1] & A[13]) , (B[1] & A[12]) , (B[1] & A[11]) , (B[1] & A[10]) , (B[1] & A[9]) ,  (B[1] & A[8]) ,  (B[1] & A[7]) ,  (B[1] & A[6]) ,  (B[1] & A[5]) ,  (B[1] & A[4]) ,  (B[1] & A[3]) ,  (B[1] & A[2]) ,  (B[1] & A[1]) ,  (B[1] & A[0]) , 1'b0 };
assign R[2][15:0] = { (B[2] & A[13]) , (B[2] & A[12]) , (B[2] & A[11]) , (B[2] & A[10]) , (B[2] & A[9]) ,  (B[2] & A[8]) ,  (B[2] & A[7]) ,  (B[2] & A[6]) ,  (B[2] & A[5]) ,  (B[2] & A[4]) ,  (B[2] & A[3]) ,  (B[2] & A[2]) ,  (B[2] & A[1]) ,  (B[2] & A[0]) , 2'b0 };
assign R[3][15:0] = { (B[3] & A[12]) , (B[3] & A[11]) , (B[3] & A[10]) , (B[3] & A[9]) ,  (B[3] & A[8]) ,  (B[3] & A[7]) ,  (B[3] & A[6]) ,  (B[3] & A[5]) ,  (B[3] & A[4]) ,  (B[3] & A[3]) ,  (B[3] & A[2]) ,  (B[3] & A[1]) ,  (B[3] & A[0]) , 3'b0 };
assign R[4][15:0] = { (B[4] & A[11]) , (B[4] & A[10]) , (B[4] & A[9]) ,  (B[4] & A[8]) ,  (B[4] & A[7]) ,  (B[4] & A[6]) ,  (B[4] & A[5]) ,  (B[4] & A[4]) ,  (B[4] & A[3]) ,  (B[4] & A[2]) ,  (B[4] & A[1]) ,  (B[4] & A[0]) , 4'b0 };
assign R[5][15:0] = { (B[5] & A[10]) , (B[5] & A[9]) ,  (B[5] & A[8]) ,  (B[5] & A[7]) ,  (B[5] & A[6]) ,  (B[5] & A[5]) ,  (B[5] & A[4]) ,  (B[5] & A[3]) ,  (B[5] & A[2]) ,  (B[5] & A[1]) ,  (B[5] & A[0]) , 5'b0 };
assign R[6][15:0] = { (B[6] & A[9]) ,  (B[6] & A[8]) ,  (B[6] & A[7]) ,  (B[6] & A[6]) ,  (B[6] & A[5]) ,  (B[6] & A[4]) ,  (B[6] & A[3]) ,  (B[6] & A[2]) ,  (B[6] & A[1]) ,  (B[6] & A[0]) , 6'b0 };
assign R[7][15:0] = { (B[7] & A[8]) ,  (B[7] & A[7]) ,  (B[7] & A[6]) ,  (B[7] & A[5]) ,  (B[7] & A[4]) ,  (B[7] & A[3]) ,  (B[7] & A[2]) ,  (B[7] & A[1]) ,  (B[7] & A[0]) , 7'b0 };
assign R[8][15:0] = { (B[8] & A[7]) ,  (B[8] & A[6]) ,  (B[8] & A[5]) ,  (B[8] & A[4]) ,  (B[8] & A[3]) ,  (B[8] & A[2]) ,  (B[8] & A[1]) ,  (B[8] & A[0]) , 8'b0 };
assign R[9][15:0] = { (B[9] & A[6]) ,  (B[9] & A[5]) ,  (B[9] & A[4]) ,  (B[9] & A[3]) ,  (B[9] & A[2]) ,  (B[9] & A[1]) ,  (B[9] & A[0]) , 9'b0 };
assign R[10][15:0] = { (B[10] & A[5]) , (B[10] & A[4]) , (B[10] & A[3]) , (B[10] & A[2]) , (B[10] & A[1]) , (B[10] & A[0]) , 10'b0 };
assign R[11][15:0] = { (B[11] & A[4]) , (B[11] & A[3]) , (B[11] & A[2]) , (B[11] & A[1]) , (B[11] & A[0]) , 11'b0 };
assign R[12][15:0] = { (B[12] & A[3]) , (B[12] & A[2]) , (B[12] & A[1]) , (B[12] & A[0]) , 12'b0 };
assign R[13][15:0] = { (B[13] & A[2]) , (B[13] & A[1]) , (B[13] & A[0]) , 13'b0 };
assign R[14][15:0] = { (B[14] & A[1]) , (B[14] & A[0]) , 14'b0 };
assign R[15][15:0] = { (B[15] & A[0]) , 15'b0 };

//assign R = R0 + R1 + R2 + R3 + R4 + R5 + R6 + R7 + R8 + R9 + R10 + R11 + R12 + R13 + R14 + R15;

endmodule