module alt_carry_look_ahead_adder_cin7
(
input [6:0] A, B,
input cin,
output [6:0] R
);
wire c0,  c1,  c2,  c3,  c4,  c5,  c6; 
wire c_one_1, c_one_2, c_one_3;
wire c_two_1, c_two_2, c_two_3, c_two_4, c_two_5, c_two_6, c_two_7;
wire c_three_1,c_three_2,c_three_3,c_three_4,c_three_5,c_three_6,c_three_7,c_three_8,c_three_9,c_three_10,c_three_11,c_three_12,c_three_13,c_three_14,c_three_15;
wire c_four_1, c_four_2, c_four_3, c_four_4, c_four_5, c_four_6, c_four_7, c_four_8, c_four_9, c_four_10, c_four_11, c_four_12, c_four_13, c_four_14, c_four_15, c_four_16, c_four_17, c_four_18, c_four_19, c_four_20, c_four_21, c_four_22, c_four_23, c_four_24, c_four_25, c_four_26, c_four_27, c_four_28, c_four_29, c_four_30, c_four_31;
wire c_five_1, c_five_2, c_five_3, c_five_4, c_five_5, c_five_6, c_five_7, c_five_8, c_five_9, c_five_10, c_five_11, c_five_12, c_five_13, c_five_14, c_five_15, c_five_16, c_five_17, c_five_18, c_five_19, c_five_20, c_five_21, c_five_22, c_five_23, c_five_24, c_five_25, c_five_26, c_five_27, c_five_28, c_five_29, c_five_30, c_five_31, c_five_32, c_five_33, c_five_34, c_five_35, c_five_36, c_five_37, c_five_38, c_five_39, c_five_40, c_five_41, c_five_42, c_five_43, c_five_44, c_five_45, c_five_46, c_five_47, c_five_48, c_five_49, c_five_50, c_five_51, c_five_52, c_five_53, c_five_54, c_five_55, c_five_56, c_five_57, c_five_58, c_five_59, c_five_60, c_five_61, c_five_62, c_five_63; 
wire c_six_1, c_six_2, c_six_3, c_six_4, c_six_5, c_six_6, c_six_7, c_six_8, c_six_9, c_six_10, c_six_11, c_six_12, c_six_13, c_six_14, c_six_15, c_six_16, c_six_17, c_six_18, c_six_19, c_six_20, c_six_21, c_six_22, c_six_23, c_six_24, c_six_25, c_six_26, c_six_27, c_six_28, c_six_29, c_six_30, c_six_31, c_six_32, c_six_33, c_six_34, c_six_35, c_six_36, c_six_37, c_six_38, c_six_39, c_six_40, c_six_41, c_six_42, c_six_43, c_six_44, c_six_45, c_six_46, c_six_47, c_six_48, c_six_49, c_six_50, c_six_51, c_six_52, c_six_53, c_six_54, c_six_55, c_six_56, c_six_57, c_six_58, c_six_59, c_six_60, c_six_61, c_six_62, c_six_63, c_six_64, c_six_65, c_six_66, c_six_67, c_six_68, c_six_69, c_six_70, c_six_71, c_six_72, c_six_73, c_six_74, c_six_75, c_six_76, c_six_77, c_six_78, c_six_79, c_six_80, c_six_81, c_six_82, c_six_83, c_six_84, c_six_85, c_six_86, c_six_87, c_six_88, c_six_89, c_six_90, c_six_91, c_six_92, c_six_93, c_six_94, c_six_95, c_six_96, c_six_97, c_six_98, c_six_99, c_six_100,  c_six_101, c_six_102, c_six_103, c_six_104, c_six_105, c_six_106, c_six_107, c_six_108, c_six_109, c_six_110, c_six_111, c_six_112, c_six_113, c_six_114, c_six_115, c_six_116, c_six_117, c_six_118, c_six_119, c_six_120, c_six_121, c_six_122, c_six_123, c_six_124, c_six_125, c_six_126, c_six_127; 



assign c0 = cin;
and(c_one_1 ,A[0],B[0]);
and(c_one_2 ,A[0],c0);
and(c_one_3 ,B[0],c0);
and(c_two_1 ,A[1],B[1]);
and(c_two_2 ,A[1],A[0],B[0]);
and(c_two_3 ,A[1],A[0],c0);
and(c_two_4 ,A[1],B[0],c0);
and(c_two_5 ,B[1],A[0],B[0]);
and(c_two_6 ,B[1],A[0],c0);
and(c_two_7 ,B[1],B[0],c0);
and(c_three_1 ,A[2],B[2]);
and(c_three_2 ,A[2],A[1],B[1]);
and(c_three_3 ,A[2],A[1],A[0],B[0]);
and(c_three_4 ,A[2],A[1],A[0],c0);
and(c_three_5 ,A[2],A[1],B[0],c0);
and(c_three_6 ,A[2],B[1],A[0],B[0]);
and(c_three_7 ,A[2],B[1],A[0],c0);
and(c_three_8 ,A[2],B[1],B[0],c0);
and(c_three_9 ,B[2],A[1],B[1]);
and(c_three_10 ,B[2],A[1],A[0],B[0]);
and(c_three_11 ,B[2],A[1],A[0],c0);
and(c_three_12 ,B[2],A[1],B[0],c0);
and(c_three_13 ,B[2],B[1],A[0],B[0]);
and(c_three_14 ,B[2],B[1],A[0],c0);
and(c_three_15 ,B[2],B[1],B[0],c0);
and(c_four_1 ,A[3],B[3]);
and(c_four_2 ,A[3],A[2],B[2]);
and(c_four_3 ,A[3],A[2],A[1],B[1]);
and(c_four_4 ,A[3],A[2],A[1],A[0],B[0]);
and(c_four_5 ,A[3],A[2],A[1],A[0],c0);
and(c_four_6 ,A[3],A[2],A[1],B[0],c0);
and(c_four_7 ,A[3],A[2],B[1],A[0],B[0]);
and(c_four_8 ,A[3],A[2],B[1],A[0],c0);
and(c_four_9 ,A[3],A[2],B[1],B[0],c0);
and(c_four_10 ,A[3],B[2],A[1],B[1]);
and(c_four_11 ,A[3],B[2],A[1],A[0],B[0]);
and(c_four_12 ,A[3],B[2],A[1],A[0],c0);
and(c_four_13 ,A[3],B[2],A[1],B[0],c0);
and(c_four_14 ,A[3],B[2],B[1],A[0],B[0]);
and(c_four_15 ,A[3],B[2],B[1],A[0],c0);
and(c_four_16 ,A[3],B[2],B[1],B[0],c0);
and(c_four_17 ,B[3],A[2],B[2]);
and(c_four_18 ,B[3],A[2],A[1],B[1]);
and(c_four_19 ,B[3],A[2],A[1],A[0],B[0]);
and(c_four_20 ,B[3],A[2],A[1],A[0],c0);
and(c_four_21 ,B[3],A[2],A[1],B[0],c0);
and(c_four_22 ,B[3],A[2],B[1],A[0],B[0]);
and(c_four_23 ,B[3],A[2],B[1],A[0],c0);
and(c_four_24 ,B[3],A[2],B[1],B[0],c0);
and(c_four_25 ,B[3],B[2],A[1],B[1]);
and(c_four_26 ,B[3],B[2],A[1],A[0],B[0]);
and(c_four_27 ,B[3],B[2],A[1],A[0],c0);
and(c_four_28 ,B[3],B[2],A[1],B[0],c0);
and(c_four_29 ,B[3],B[2],B[1],A[0],B[0]);
and(c_four_30 ,B[3],B[2],B[1],A[0],c0);
and(c_four_31 ,B[3],B[2],B[1],B[0],c0);
and(c_five_1 ,A[4],B[4]);
and(c_five_2 ,A[4],A[3],B[3]);
and(c_five_3 ,A[4],A[3],A[2],B[2]);
and(c_five_4 ,A[4],A[3],A[2],A[1],B[1]);
and(c_five_5 ,A[4],A[3],A[2],A[1],A[0],B[0]);
and(c_five_6 ,A[4],A[3],A[2],A[1],A[0],c0);
and(c_five_7 ,A[4],A[3],A[2],A[1],B[0],c0);
and(c_five_8 ,A[4],A[3],A[2],B[1],A[0],B[0]);
and(c_five_9 ,A[4],A[3],A[2],B[1],A[0],c0);
and(c_five_10 ,A[4],A[3],A[2],B[1],B[0],c0);
and(c_five_11 ,A[4],A[3],B[2],A[1],B[1]);
and(c_five_12 ,A[4],A[3],B[2],A[1],A[0],B[0]);
and(c_five_13 ,A[4],A[3],B[2],A[1],A[0],c0);
and(c_five_14 ,A[4],A[3],B[2],A[1],B[0],c0);
and(c_five_15 ,A[4],A[3],B[2],B[1],A[0],B[0]);
and(c_five_16 ,A[4],A[3],B[2],B[1],A[0],c0);
and(c_five_17 ,A[4],A[3],B[2],B[1],B[0],c0);
and(c_five_18 ,A[4],B[3],A[2],B[2]);
and(c_five_19 ,A[4],B[3],A[2],A[1],B[1]);
and(c_five_20 ,A[4],B[3],A[2],A[1],A[0],B[0]);
and(c_five_21 ,A[4],B[3],A[2],A[1],A[0],c0);
and(c_five_22 ,A[4],B[3],A[2],A[1],B[0],c0);
and(c_five_23 ,A[4],B[3],A[2],B[1],A[0],B[0]);
and(c_five_24 ,A[4],B[3],A[2],B[1],A[0],c0);
and(c_five_25 ,A[4],B[3],A[2],B[1],B[0],c0);
and(c_five_26 ,A[4],B[3],B[2],A[1],B[1]);
and(c_five_27 ,A[4],B[3],B[2],A[1],A[0],B[0]);
and(c_five_28 ,A[4],B[3],B[2],A[1],A[0],c0);
and(c_five_29 ,A[4],B[3],B[2],A[1],B[0],c0);
and(c_five_30 ,A[4],B[3],B[2],B[1],A[0],B[0]);
and(c_five_31 ,A[4],B[3],B[2],B[1],A[0],c0);
and(c_five_32 ,A[4],B[3],B[2],B[1],B[0],c0);
and(c_five_33 ,B[4],A[3],B[3]);
and(c_five_34 ,B[4],A[3],A[2],B[2]);
and(c_five_35 ,B[4],A[3],A[2],A[1],B[1]);
and(c_five_36 ,B[4],A[3],A[2],A[1],A[0],B[0]);
and(c_five_37 ,B[4],A[3],A[2],A[1],A[0],c0);
and(c_five_38 ,B[4],A[3],A[2],A[1],B[0],c0);
and(c_five_39 ,B[4],A[3],A[2],B[1],A[0],B[0]);
and(c_five_40 ,B[4],A[3],A[2],B[1],A[0],c0);
and(c_five_41 ,B[4],A[3],A[2],B[1],B[0],c0);
and(c_five_42 ,B[4],A[3],B[2],A[1],B[1]);
and(c_five_43 ,B[4],A[3],B[2],A[1],A[0],B[0]);
and(c_five_44 ,B[4],A[3],B[2],A[1],A[0],c0);
and(c_five_45 ,B[4],A[3],B[2],A[1],B[0],c0);
and(c_five_46 ,B[4],A[3],B[2],B[1],A[0],B[0]);
and(c_five_47 ,B[4],A[3],B[2],B[1],A[0],c0);
and(c_five_48 ,B[4],A[3],B[2],B[1],B[0],c0);
and(c_five_49 ,B[4],B[3],A[2],B[2]);
and(c_five_50 ,B[4],B[3],A[2],A[1],B[1]);
and(c_five_51 ,B[4],B[3],A[2],A[1],A[0],B[0]);
and(c_five_52 ,B[4],B[3],A[2],A[1],A[0],c0);
and(c_five_53 ,B[4],B[3],A[2],A[1],B[0],c0);
and(c_five_54 ,B[4],B[3],A[2],B[1],A[0],B[0]);
and(c_five_55 ,B[4],B[3],A[2],B[1],A[0],c0);
and(c_five_56 ,B[4],B[3],A[2],B[1],B[0],c0);
and(c_five_57 ,B[4],B[3],B[2],A[1],B[1]);
and(c_five_58 ,B[4],B[3],B[2],A[1],A[0],B[0]);
and(c_five_59 ,B[4],B[3],B[2],A[1],A[0],c0);
and(c_five_60 ,B[4],B[3],B[2],A[1],B[0],c0);
and(c_five_61 ,B[4],B[3],B[2],B[1],A[0],B[0]);
and(c_five_62 ,B[4],B[3],B[2],B[1],A[0],c0);
and(c_five_63 ,B[4],B[3],B[2],B[1],B[0],c0);
and(c_six_1 ,A[5],B[5]);
and(c_six_2 ,A[5],A[4],B[4]);
and(c_six_3 ,A[5],A[4],A[3],B[3]);
and(c_six_4 ,A[5],A[4],A[3],A[2],B[2]);
and(c_six_5 ,A[5],A[4],A[3],A[2],A[1],B[1]);
and(c_six_6 ,A[5],A[4],A[3],A[2],A[1],A[0],B[0]);
and(c_six_7 ,A[5],A[4],A[3],A[2],A[1],A[0],c0);
and(c_six_8 ,A[5],A[4],A[3],A[2],A[1],B[0],c0);
and(c_six_9 ,A[5],A[4],A[3],A[2],B[1],A[0],B[0]);
and(c_six_10 ,A[5],A[4],A[3],A[2],B[1],A[0],c0);
and(c_six_11 ,A[5],A[4],A[3],A[2],B[1],B[0],c0);
and(c_six_12 ,A[5],A[4],A[3],B[2],A[1],B[1]);
and(c_six_13 ,A[5],A[4],A[3],B[2],A[1],A[0],B[0]);
and(c_six_14 ,A[5],A[4],A[3],B[2],A[1],A[0],c0);
and(c_six_15 ,A[5],A[4],A[3],B[2],A[1],B[0],c0);
and(c_six_16 ,A[5],A[4],A[3],B[2],B[1],A[0],B[0]);
and(c_six_17 ,A[5],A[4],A[3],B[2],B[1],A[0],c0);
and(c_six_18 ,A[5],A[4],A[3],B[2],B[1],B[0],c0);
and(c_six_19 ,A[5],A[4],B[3],A[2],B[2]);
and(c_six_20 ,A[5],A[4],B[3],A[2],A[1],B[1]);
and(c_six_21 ,A[5],A[4],B[3],A[2],A[1],A[0],B[0]);
and(c_six_22 ,A[5],A[4],B[3],A[2],A[1],A[0],c0);
and(c_six_23 ,A[5],A[4],B[3],A[2],A[1],B[0],c0);
and(c_six_24 ,A[5],A[4],B[3],A[2],B[1],A[0],B[0]);
and(c_six_25 ,A[5],A[4],B[3],A[2],B[1],A[0],c0);
and(c_six_26 ,A[5],A[4],B[3],A[2],B[1],B[0],c0);
and(c_six_27 ,A[5],A[4],B[3],B[2],A[1],B[1]);
and(c_six_28 ,A[5],A[4],B[3],B[2],A[1],A[0],B[0]);
and(c_six_29 ,A[5],A[4],B[3],B[2],A[1],A[0],c0);
and(c_six_30 ,A[5],A[4],B[3],B[2],A[1],B[0],c0);
and(c_six_31 ,A[5],A[4],B[3],B[2],B[1],A[0],B[0]);
and(c_six_32 ,A[5],A[4],B[3],B[2],B[1],A[0],c0);
and(c_six_33 ,A[5],A[4],B[3],B[2],B[1],B[0],c0);
and(c_six_34 ,A[5],B[4],A[3],B[3]);
and(c_six_35 ,A[5],B[4],A[3],A[2],B[2]);
and(c_six_36 ,A[5],B[4],A[3],A[2],A[1],B[1]);
and(c_six_37 ,A[5],B[4],A[3],A[2],A[1],A[0],B[0]);
and(c_six_38 ,A[5],B[4],A[3],A[2],A[1],A[0],c0);
and(c_six_39 ,A[5],B[4],A[3],A[2],A[1],B[0],c0);
and(c_six_40 ,A[5],B[4],A[3],A[2],B[1],A[0],B[0]);
and(c_six_41 ,A[5],B[4],A[3],A[2],B[1],A[0],c0);
and(c_six_42 ,A[5],B[4],A[3],A[2],B[1],B[0],c0);
and(c_six_43 ,A[5],B[4],A[3],B[2],A[1],B[1]);
and(c_six_44 ,A[5],B[4],A[3],B[2],A[1],A[0],B[0]);
and(c_six_45 ,A[5],B[4],A[3],B[2],A[1],A[0],c0);
and(c_six_46 ,A[5],B[4],A[3],B[2],A[1],B[0],c0);
and(c_six_47 ,A[5],B[4],A[3],B[2],B[1],A[0],B[0]);
and(c_six_48 ,A[5],B[4],A[3],B[2],B[1],A[0],c0);
and(c_six_49 ,A[5],B[4],A[3],B[2],B[1],B[0],c0);
and(c_six_50 ,A[5],B[4],B[3],A[2],B[2]);
and(c_six_51 ,A[5],B[4],B[3],A[2],A[1],B[1]);
and(c_six_52 ,A[5],B[4],B[3],A[2],A[1],A[0],B[0]);
and(c_six_53 ,A[5],B[4],B[3],A[2],A[1],A[0],c0);
and(c_six_54 ,A[5],B[4],B[3],A[2],A[1],B[0],c0);
and(c_six_55 ,A[5],B[4],B[3],A[2],B[1],A[0],B[0]);
and(c_six_56 ,A[5],B[4],B[3],A[2],B[1],A[0],c0);
and(c_six_57 ,A[5],B[4],B[3],A[2],B[1],B[0],c0);
and(c_six_58 ,A[5],B[4],B[3],B[2],A[1],B[1]);
and(c_six_59 ,A[5],B[4],B[3],B[2],A[1],A[0],B[0]);
and(c_six_60 ,A[5],B[4],B[3],B[2],A[1],A[0],c0);
and(c_six_61 ,A[5],B[4],B[3],B[2],A[1],B[0],c0);
and(c_six_62 ,A[5],B[4],B[3],B[2],B[1],A[0],B[0]);
and(c_six_63 ,A[5],B[4],B[3],B[2],B[1],A[0],c0);
and(c_six_64 ,A[5],B[4],B[3],B[2],B[1],B[0],c0);
and(c_six_65 ,B[5],A[4],B[4]);
and(c_six_66 ,B[5],A[4],A[3],B[3]);
and(c_six_67 ,B[5],A[4],A[3],A[2],B[2]);
and(c_six_68 ,B[5],A[4],A[3],A[2],A[1],B[1]);
and(c_six_69 ,B[5],A[4],A[3],A[2],A[1],A[0],B[0]);
and(c_six_70 ,B[5],A[4],A[3],A[2],A[1],A[0],c0);
and(c_six_71 ,B[5],A[4],A[3],A[2],A[1],B[0],c0);
and(c_six_72 ,B[5],A[4],A[3],A[2],B[1],A[0],B[0]);
and(c_six_73 ,B[5],A[4],A[3],A[2],B[1],A[0],c0);
and(c_six_74 ,B[5],A[4],A[3],A[2],B[1],B[0],c0);
and(c_six_75 ,B[5],A[4],A[3],B[2],A[1],B[1]);
and(c_six_76 ,B[5],A[4],A[3],B[2],A[1],A[0],B[0]);
and(c_six_77 ,B[5],A[4],A[3],B[2],A[1],A[0],c0);
and(c_six_78 ,B[5],A[4],A[3],B[2],A[1],B[0],c0);
and(c_six_79 ,B[5],A[4],A[3],B[2],B[1],A[0],B[0]);
and(c_six_80 ,B[5],A[4],A[3],B[2],B[1],A[0],c0);
and(c_six_81 ,B[5],A[4],A[3],B[2],B[1],B[0],c0);
and(c_six_82 ,B[5],A[4],B[3],A[2],B[2]);
and(c_six_83 ,B[5],A[4],B[3],A[2],A[1],B[1]);
and(c_six_84 ,B[5],A[4],B[3],A[2],A[1],A[0],B[0]);
and(c_six_85 ,B[5],A[4],B[3],A[2],A[1],A[0],c0);
and(c_six_86 ,B[5],A[4],B[3],A[2],A[1],B[0],c0);
and(c_six_87 ,B[5],A[4],B[3],A[2],B[1],A[0],B[0]);
and(c_six_88 ,B[5],A[4],B[3],A[2],B[1],A[0],c0);
and(c_six_89 ,B[5],A[4],B[3],A[2],B[1],B[0],c0);
and(c_six_90 ,B[5],A[4],B[3],B[2],A[1],B[1]);
and(c_six_91 ,B[5],A[4],B[3],B[2],A[1],A[0],B[0]);
and(c_six_92 ,B[5],A[4],B[3],B[2],A[1],A[0],c0);
and(c_six_93 ,B[5],A[4],B[3],B[2],A[1],B[0],c0);
and(c_six_94 ,B[5],A[4],B[3],B[2],B[1],A[0],B[0]);
and(c_six_95 ,B[5],A[4],B[3],B[2],B[1],A[0],c0);
and(c_six_96 ,B[5],A[4],B[3],B[2],B[1],B[0],c0);
and(c_six_97 ,B[5],B[4],A[3],B[3]);
and(c_six_98 ,B[5],B[4],A[3],A[2],B[2]);
and(c_six_99 ,B[5],B[4],A[3],A[2],A[1],B[1]);
and(c_six_100 ,B[5],B[4],A[3],A[2],A[1],A[0],B[0]);
and(c_six_101 ,B[5],B[4],A[3],A[2],A[1],A[0],c0);
and(c_six_102 ,B[5],B[4],A[3],A[2],A[1],B[0],c0);
and(c_six_103 ,B[5],B[4],A[3],A[2],B[1],A[0],B[0]);
and(c_six_104 ,B[5],B[4],A[3],A[2],B[1],A[0],c0);
and(c_six_105 ,B[5],B[4],A[3],A[2],B[1],B[0],c0);
and(c_six_106 ,B[5],B[4],A[3],B[2],A[1],B[1]);
and(c_six_107 ,B[5],B[4],A[3],B[2],A[1],A[0],B[0]);
and(c_six_108 ,B[5],B[4],A[3],B[2],A[1],A[0],c0);
and(c_six_109 ,B[5],B[4],A[3],B[2],A[1],B[0],c0);
and(c_six_110 ,B[5],B[4],A[3],B[2],B[1],A[0],B[0]);
and(c_six_111 ,B[5],B[4],A[3],B[2],B[1],A[0],c0);
and(c_six_112 ,B[5],B[4],A[3],B[2],B[1],B[0],c0);
and(c_six_113 ,B[5],B[4],B[3],A[2],B[2]);
and(c_six_114 ,B[5],B[4],B[3],A[2],A[1],B[1]);
and(c_six_115 ,B[5],B[4],B[3],A[2],A[1],A[0],B[0]);
and(c_six_116 ,B[5],B[4],B[3],A[2],A[1],A[0],c0);
and(c_six_117 ,B[5],B[4],B[3],A[2],A[1],B[0],c0);
and(c_six_118 ,B[5],B[4],B[3],A[2],B[1],A[0],B[0]);
and(c_six_119 ,B[5],B[4],B[3],A[2],B[1],A[0],c0);
and(c_six_120 ,B[5],B[4],B[3],A[2],B[1],B[0],c0);
and(c_six_121 ,B[5],B[4],B[3],B[2],A[1],B[1]);
and(c_six_122 ,B[5],B[4],B[3],B[2],A[1],A[0],B[0]);
and(c_six_123 ,B[5],B[4],B[3],B[2],A[1],A[0],c0);
and(c_six_124 ,B[5],B[4],B[3],B[2],A[1],B[0],c0);
and(c_six_125 ,B[5],B[4],B[3],B[2],B[1],A[0],B[0]);
and(c_six_126 ,B[5],B[4],B[3],B[2],B[1],A[0],c0);
and(c_six_127 ,B[5],B[4],B[3],B[2],B[1],B[0],c0);




assign c1 = c_one_1| c_one_2| c_one_3;
assign c2 = c_two_1| c_two_2| c_two_3| c_two_4| c_two_5| c_two_6| c_two_7;
assign c3 = c_three_1|c_three_2|c_three_3|c_three_4|c_three_5|c_three_6|c_three_7|c_three_8|c_three_9|c_three_10|c_three_11|c_three_12|c_three_13|c_three_14|c_three_15;
assign c4 = c_four_1| c_four_2| c_four_3| c_four_4| c_four_5| c_four_6| c_four_7| c_four_8| c_four_9| c_four_10| c_four_11| c_four_12| c_four_13| c_four_14| c_four_15| c_four_16| c_four_17| c_four_18| c_four_19| c_four_20| c_four_21| c_four_22| c_four_23| c_four_24| c_four_25| c_four_26| c_four_27| c_four_28| c_four_29| c_four_30| c_four_31;
assign c5 = c_five_1| c_five_2| c_five_3| c_five_4| c_five_5| c_five_6| c_five_7| c_five_8| c_five_9| c_five_10| c_five_11| c_five_12| c_five_13| c_five_14| c_five_15| c_five_16| c_five_17| c_five_18| c_five_19| c_five_20| c_five_21| c_five_22| c_five_23| c_five_24| c_five_25| c_five_26| c_five_27| c_five_28| c_five_29| c_five_30| c_five_31| c_five_32| c_five_33| c_five_34| c_five_35| c_five_36| c_five_37| c_five_38| c_five_39| c_five_40| c_five_41| c_five_42| c_five_43| c_five_44| c_five_45| c_five_46| c_five_47| c_five_48| c_five_49| c_five_50| c_five_51| c_five_52| c_five_53| c_five_54| c_five_55| c_five_56| c_five_57| c_five_58| c_five_59| c_five_60| c_five_61| c_five_62| c_five_63; 
assign c6 = c_six_1| c_six_2| c_six_3| c_six_4| c_six_5| c_six_6| c_six_7| c_six_8| c_six_9| c_six_10| c_six_11| c_six_12| c_six_13| c_six_14| c_six_15| c_six_16| c_six_17| c_six_18| c_six_19| c_six_20| c_six_21| c_six_22| c_six_23| c_six_24| c_six_25| c_six_26| c_six_27| c_six_28| c_six_29| c_six_30| c_six_31| c_six_32| c_six_33| c_six_34| c_six_35| c_six_36| c_six_37| c_six_38| c_six_39| c_six_40| c_six_41| c_six_42| c_six_43| c_six_44| c_six_45| c_six_46| c_six_47| c_six_48| c_six_49| c_six_50| c_six_51| c_six_52| c_six_53| c_six_54| c_six_55| c_six_56| c_six_57| c_six_58| c_six_59| c_six_60| c_six_61| c_six_62| c_six_63| c_six_64| c_six_65| c_six_66| c_six_67| c_six_68| c_six_69| c_six_70| c_six_71| c_six_72| c_six_73| c_six_74| c_six_75| c_six_76| c_six_77| c_six_78| c_six_79| c_six_80| c_six_81| c_six_82| c_six_83| c_six_84| c_six_85| c_six_86| c_six_87| c_six_88| c_six_89| c_six_90| c_six_91| c_six_92| c_six_93| c_six_94| c_six_95| c_six_96| c_six_97| c_six_98| c_six_99| c_six_100|  c_six_101| c_six_102| c_six_103| c_six_104| c_six_105| c_six_106| c_six_107| c_six_108| c_six_109| c_six_110| c_six_111| c_six_112| c_six_113| c_six_114| c_six_115| c_six_116| c_six_117| c_six_118| c_six_119| c_six_120| c_six_121| c_six_122| c_six_123| c_six_124| c_six_125| c_six_126| c_six_127; 






assign R[0] = A[0] ^ B[0] ^ c0;
assign R[1] = A[1] ^ B[1] ^ c1;
assign R[2] = A[2] ^ B[2] ^ c2;
assign R[3] = A[3] ^ B[3] ^ c3;
assign R[4] = A[4] ^ B[4] ^ c4;
assign R[5] = A[5] ^ B[5] ^ c5;
assign R[6] = A[6] ^ B[6] ^ c6;


endmodule
