module simple16adder
(
input [15:0] A, B,
output [15:0] res
);

assign res = A + B;

endmodule