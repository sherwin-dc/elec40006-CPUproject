module alt_carry_look_ahead_adder_cin
(
input [15:0] A, B,
input cin,
output [15:0] R
);
wire p0,  p1,  p2,  p3,  p4,  p5,  p6,  p7,  p8,  p9,  p10, p11, p12, p13, p14, p15; 
wire c0,  c1,  c2,  c3,  c4,  c5,  c6,  c7,  c8,  c9,  c10, c11, c12, c13, c14, c15; 
wire [15:0] c_fiften;
wire [14:0] c_fourtn;
wire [13:0] c_thirtn;
wire [12:0] c_twelve;
wire [11:0] c_eleven;
wire [10:0] c_ten;
wire [9:0] c_nine;
wire [8:0] c_eight;
wire [7:0] c_seven;
wire [6:0] c_six;
wire [5:0] c_five;
wire [4:0] c_four;
wire [3:0] c_three;
wire [2:0] c_two;
wire [1:0] c_one;

assign p0 = A[0] ^ B[0];
assign p1 = A[1] ^ B[1];
assign p2 = A[2] ^ B[2];
assign p3 = A[3] ^ B[3];
assign p4 = A[4] ^ B[4];
assign p5 = A[5] ^ B[5];
assign p6 = A[6] ^ B[6];
assign p7 = A[7] ^ B[7];
assign p8 = A[8] ^ B[8];
assign p9 = A[9] ^ B[9];
assign p10 = A[10] ^ B[10];
assign p11 = A[11] ^ B[11];
assign p12 = A[12] ^ B[12];
assign p13 = A[13] ^ B[13];
assign p14 = A[14] ^ B[14];
assign p15 = A[15] ^ B[15];


assign c0 = cin;
and(c_one[0] , A[0] , B[0]); 
 and(c_one[1] , p0 , cin);
and(c_two[0] , A[1] , B[1]); 
 and(c_two[1] , p1 , A[0] , B[0]); 
 and(c_two[2] , p1 , p0 , cin);
and(c_three[0] , A[2] , B[2]); 
 and(c_three[1] , p2 , A[1] , B[1]); 
 and(c_three[2] , p2 , p1 , A[0] , B[0]); 
 and(c_three[3] , p2 , p1 , p0 , cin);
and(c_four[0] , A[3] , B[3]); 
 and(c_four[1] , p3 , A[2] , B[2]); 
 and(c_four[2] , p3 , p2 , A[1] , B[1]); 
 and(c_four[3] , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_four[4] , p3 , p2 , p1 , p0 , cin);
and(c_five[0] , A[4] , B[4]); 
 and(c_five[1] , p4 , A[3] , B[3]); 
 and(c_five[2] , p4 , p3 , A[2] , B[2]); 
 and(c_five[3] , p4 , p3 , p2 , A[1] , B[1]); 
 and(c_five[4] , p4 , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_five[5] , p4 , p3 , p2 , p1 , p0 , cin);
and(c_six[0] , A[5] , B[5]); 
 and(c_six[1] , p5 , A[4] , B[4]); 
 and(c_six[2] , p5 , p4 , A[3] , B[3]); 
 and(c_six[3] , p5 , p4 , p3 , A[2] , B[2]); 
 and(c_six[4] , p5 , p4 , p3 , p2 , A[1] , B[1]); 
 and(c_six[5] , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_six[6] , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_seven[0] , A[6] , B[6]); 
 and(c_seven[1] , p6 , A[5] , B[5]); 
 and(c_seven[2] , p6 , p5 , A[4] , B[4]); 
 and(c_seven[3] , p6 , p5 , p4 , A[3] , B[3]); 
 and(c_seven[4] , p6 , p5 , p4 , p3 , A[2] , B[2]); 
 and(c_seven[5] , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
 and(c_seven[6] , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_seven[7] , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_eight[0] , A[7] , B[7]); 
 and(c_eight[1] , p7 , A[6] , B[6]); 
 and(c_eight[2] , p7 , p6 , A[5] , B[5]); 
 and(c_eight[3] , p7 , p6 , p5 , A[4] , B[4]); 
 and(c_eight[4] , p7 , p6 , p5 , p4 , A[3] , B[3]); 
 and(c_eight[5] , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
 and(c_eight[6] , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
 and(c_eight[7] , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_eight[8] , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_nine[0] , A[8] , B[8]); 
 and(c_nine[1] , p8 , A[7] , B[7]); 
 and(c_nine[2] , p8 , p7 , A[6] , B[6]); 
 and(c_nine[3] , p8 , p7 , p6 , A[5] , B[5]); 
 and(c_nine[4] , p8 , p7 , p6 , p5 , A[4] , B[4]); 
 and(c_nine[5] , p8 , p7 , p6 , p5 , p4 , A[3] , B[3]); 
 and(c_nine[6] , p8 , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
 and(c_nine[7] , p8 , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
 and(c_nine[8] , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_nine[9] , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_ten[0] , A[9] , B[9]); 
 and(c_ten[1] , p9 , A[8] , B[8]); 
 and(c_ten[2] , p9 , p8 , A[7] , B[7]); 
 and(c_ten[3] , p9 , p8 , p7 , A[6] , B[6]); 
 and(c_ten[4] , p9 , p8 , p7 , p6 , A[5] , B[5]); 
 and(c_ten[5] , p9 , p8 , p7 , p6 , p5 , A[4] , B[4]); 
 and(c_ten[6] , p9 , p8 , p7 , p6 , p5 , p4 , A[3] , B[3]); 
 and(c_ten[7] , p9 , p8 , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
 and(c_ten[8] , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
 and(c_ten[9] , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_ten[10] , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_eleven[0] , A[10] , B[10]); 
 and(c_eleven[1] , p10 , A[9] , B[9]); 
 and(c_eleven[2] , p10 , p9 , A[8] , B[8]); 
 and(c_eleven[3] , p10 , p9 , p8 , A[7] , B[7]); 
 and(c_eleven[4] , p10 , p9 , p8 , p7 , A[6] , B[6]); 
 and(c_eleven[5] , p10 , p9 , p8 , p7 , p6 , A[5] , B[5]); 
 and(c_eleven[6] , p10 , p9 , p8 , p7 , p6 , p5 , A[4] , B[4]); 
 and(c_eleven[7] , p10 , p9 , p8 , p7 , p6 , p5 , p4 , A[3] , B[3]); 
 and(c_eleven[8] , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
 and(c_eleven[9] , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
 and(c_eleven[10] , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
 and(c_eleven[11] , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_twelve[0] , A[11] , B[11]); 
and(c_twelve[1] , p11 , A[10] , B[10]); 
and(c_twelve[2] , p11 , p10 , A[9] , B[9]); 
and(c_twelve[3] , p11 , p10 , p9 , A[8] , B[8]); 
and(c_twelve[4] , p11 , p10 , p9 , p8 , A[7] , B[7]); 
and(c_twelve[5] , p11 , p10 , p9 , p8 , p7 , A[6] , B[6]); 
and(c_twelve[6] , p11 , p10 , p9 , p8 , p7 , p6 , A[5] , B[5]); 
and(c_twelve[7] , p11 , p10 , p9 , p8 , p7 , p6 , p5 , A[4] , B[4]); 
and(c_twelve[8] , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , A[3] , B[3]); 
and(c_twelve[9] , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
and(c_twelve[10] , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
and(c_twelve[11] ,p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
and(c_twelve[12] ,p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_thirtn[0] , A[12] , B[12]); 
and(c_thirtn[1] , p12 , A[11] , B[11]); 
and(c_thirtn[2] , p12 , p11 , A[10] , B[10]); 
and(c_thirtn[3] , p12 , p11 , p10 , A[9] , B[9]); 
and(c_thirtn[4] , p12 , p11 , p10 , p9 , A[8] , B[8]); 
and(c_thirtn[5] , p12 , p11 , p10 , p9 , p8 , A[7] , B[7]); 
and(c_thirtn[6] , p12 , p11 , p10 , p9 , p8 , p7 , A[6] , B[6]); 
and(c_thirtn[7] , p12 , p11 , p10 , p9 , p8 , p7 , p6 , A[5] , B[5]); 
and(c_thirtn[8] , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , A[4] , B[4]); 
and(c_thirtn[9] , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , A[3] , B[3]); 
and(c_thirtn[10] , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
and(c_thirtn[11] ,p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
and(c_thirtn[12] ,p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
and(c_thirtn[13] ,p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_fourtn[0] , A[13] , B[13]); 
and(c_fourtn[1] , p13 , A[12] , B[12]); 
and(c_fourtn[2] , p13 , p12 , A[11] , B[11]); 
and(c_fourtn[3] , p13 , p12 , p11 , A[10] , B[10]); 
and(c_fourtn[4] , p13 , p12 , p11 , p10 , A[9] , B[9]); 
and(c_fourtn[5] , p13 , p12 , p11 , p10 , p9 , A[8] , B[8]); 
and(c_fourtn[6] , p13 , p12 , p11 , p10 , p9 , p8 , A[7] , B[7]); 
and(c_fourtn[7] , p13 , p12 , p11 , p10 , p9 , p8 , p7 , A[6] , B[6]); 
and(c_fourtn[8] , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , A[5] , B[5]); 
and(c_fourtn[9] , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , A[4] , B[4]); 
and(c_fourtn[10] , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , A[3] , B[3]); 
and(c_fourtn[11] ,p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
and(c_fourtn[12] ,p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
and(c_fourtn[13] ,p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
and(c_fourtn[14] ,p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);
and(c_fiften[0] , A[14] , B[14]); 
and(c_fiften[1] , p14 , A[13] , B[13]); 
and(c_fiften[2] , p14 , p13 , A[12] , B[12]); 
and(c_fiften[3] , p14 , p13 , p12 , A[11] , B[11]); 
and(c_fiften[4] , p14 , p13 , p12 , p11 , A[10] , B[10]); 
and(c_fiften[5] , p14 , p13 , p12 , p11 , p10 , A[9] , B[9]); 
and(c_fiften[6] , p14 , p13 , p12 , p11 , p10 , p9 , A[8] , B[8]); 
and(c_fiften[7] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , A[7] , B[7]); 
and(c_fiften[8] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , A[6] , B[6]); 
and(c_fiften[9] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , A[5] , B[5]); 
and(c_fiften[10] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , A[4] , B[4]); 
and(c_fiften[11] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , A[3] , B[3]); 
and(c_fiften[12] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , A[2] , B[2]); 
and(c_fiften[13] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , A[1] , B[1]); 
and(c_fiften[14] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , A[0] , B[0]); 
and(c_fiften[15] , p14 , p13 , p12 , p11 , p10 , p9 , p8 , p7 , p6 , p5 , p4 , p3 , p2 , p1 , p0 , cin);

assign c1 = c_one[0] | c_one[1];
assign c2 = c_two[0] | c_two[1] | c_two[2]; 
assign c3 = c_three[0] | c_three[1] | c_three[2] | c_three[3]; 
assign c4 = c_four[0] | c_four[1] | c_four[2] | c_four[3] | c_four[4];
assign c5 = c_five[0] | c_five[1] | c_five[2] | c_five[3] | c_five[4] | c_five[5];
assign c6 = c_six[0] | c_six[1] | c_six[2] | c_six[3] | c_six[4] | c_six[5] | c_six[6];
assign c7 = c_seven[0] | c_seven[1] | c_seven[2] | c_seven[3] | c_seven[4] | c_seven[5] | c_seven[6] | c_seven[7]; 
assign c8 = c_eight[0] | c_eight[1] | c_eight[2] | c_eight[3] | c_eight[4] | c_eight[5] | c_eight[6] | c_eight[7] | c_eight[8];
assign c9 = c_nine[0] | c_nine[1] | c_nine[2] | c_nine[3] | c_nine[4] | c_nine[5] | c_nine[6] | c_nine[7] | c_nine[8] | c_nine[9]; 
assign c10 = c_ten[0] | c_ten[1] | c_ten[2] | c_ten[3] | c_ten[4] | c_ten[5] | c_ten[6] | c_ten[7] | c_ten[8] | c_ten[9] | c_ten[10];
assign c11 = c_eleven[0] | c_eleven[1] | c_eleven[2] | c_eleven[3] | c_eleven[4] | c_eleven[5] | c_eleven[6] | c_eleven[7] | c_eleven[8] | c_eleven[9] | c_eleven[10] | c_eleven[11];
assign c12 = c_twelve[0] | c_twelve[1] | c_twelve[2] | c_twelve[3] | c_twelve[4] | c_twelve[5] | c_twelve[6] | c_twelve[7] | c_twelve[8] | c_twelve[9] | c_twelve[10] | c_twelve[11] | c_twelve[12];
assign c13 = c_thirtn[0] | c_thirtn[1] | c_thirtn[2] | c_thirtn[3] | c_thirtn[4] | c_thirtn[5] | c_thirtn[6] | c_thirtn[7] | c_thirtn[8] | c_thirtn[9] | c_thirtn[10] | c_thirtn[11] | c_thirtn[12] | c_thirtn[13];
assign c14 = c_fourtn[0] | c_fourtn[1] | c_fourtn[2] | c_fourtn[3] | c_fourtn[4] | c_fourtn[5] | c_fourtn[6] | c_fourtn[7] | c_fourtn[8] | c_fourtn[9] | c_fourtn[10] |c_fourtn[11] |c_fourtn[12] |c_fourtn[13] |c_fourtn[14];
assign c15 = c_fiften[0] | c_fiften[1] | c_fiften[2] | c_fiften[3] | c_fiften[4] | c_fiften[5] | c_fiften[6] | c_fiften[7] | c_fiften[8] | c_fiften[9] | c_fiften[10] | c_fiften[11] | c_fiften[12] | c_fiften[13] | c_fiften[14] | c_fiften[15];

assign R[0] = p0 ^ c0;
assign R[1] = p1 ^ c1;
assign R[2] = p2 ^ c2;
assign R[3] = p3 ^ c3;
assign R[4] = p4 ^ c4;
assign R[5] = p5 ^ c5;
assign R[6] = p6 ^ c6;
assign R[7] = p7 ^ c7;
assign R[8] = p8 ^ c8;
assign R[9] = p9 ^ c9;
assign R[10] = p10 ^ c10;
assign R[11] = p11 ^ c11;
assign R[12] = p12 ^ c12;
assign R[13] = p13 ^ c13;
assign R[14] = p14 ^ c14;
assign R[15] = p15 ^ c15;

endmodule