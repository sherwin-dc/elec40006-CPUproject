module two_CLA8_adders
(

input [15:0] A, B,
input cin
);
endmodule
