module new_carry_look_ahead_adder_cin7
(
input [6:0] A, B,
input cin,
output [6:0] R
);
wire c0,  c1,  c2,  c3,  c4,  c5,  c6; 





assign c0 = cin;
assign c1 = (A[0]&B[0])|(A[0]&c0)|(B[0]&c0);
assign c2 = (A[1]&B[1])|(A[1]&A[0]&B[0])|(A[1]&A[0]&c0)|(A[1]&B[0]&c0)|(B[1]&A[0]&B[0])|(B[1]&A[0]&c0)|(B[1]&B[0]&c0);
assign c3 = (A[2]&B[2])|(A[2]&A[1]&B[1])|(A[2]&A[1]&A[0]&B[0])|(A[2]&A[1]&A[0]&c0)|(A[2]&A[1]&B[0]&c0)|(A[2]&B[1]&A[0]&B[0])|(A[2]&B[1]&A[0]&c0)|(A[2]&B[1]&B[0]&c0)|(B[2]&A[1]&B[1])|(B[2]&A[1]&A[0]&B[0])|(B[2]&A[1]&A[0]&c0)|(B[2]&A[1]&B[0]&c0)|(B[2]&B[1]&A[0]&B[0])|(B[2]&B[1]&A[0]&c0)|(B[2]&B[1]&B[0]&c0);
assign c4 = (A[3]&B[3])|(A[3]&A[2]&B[2])|(A[3]&A[2]&A[1]&B[1])|(A[3]&A[2]&A[1]&A[0]&B[0])|(A[3]&A[2]&A[1]&A[0]&c0)|(A[3]&A[2]&A[1]&B[0]&c0)|(A[3]&A[2]&B[1]&A[0]&B[0])|(A[3]&A[2]&B[1]&A[0]&c0)|(A[3]&A[2]&B[1]&B[0]&c0)|(A[3]&B[2]&A[1]&B[1])|(A[3]&B[2]&A[1]&A[0]&B[0])|(A[3]&B[2]&A[1]&A[0]&c0)|(A[3]&B[2]&A[1]&B[0]&c0)|(A[3]&B[2]&B[1]&A[0]&B[0])|(A[3]&B[2]&B[1]&A[0]&c0)|(A[3]&B[2]&B[1]&B[0]&c0)|(B[3]&A[2]&B[2])|(B[3]&A[2]&A[1]&B[1])|(B[3]&A[2]&A[1]&A[0]&B[0])|(B[3]&A[2]&A[1]&A[0]&c0)|(B[3]&A[2]&A[1]&B[0]&c0)|(B[3]&A[2]&B[1]&A[0]&B[0])|(B[3]&A[2]&B[1]&A[0]&c0)|(B[3]&A[2]&B[1]&B[0]&c0)|(B[3]&B[2]&A[1]&B[1])|(B[3]&B[2]&A[1]&A[0]&B[0])|(B[3]&B[2]&A[1]&A[0]&c0)|(B[3]&B[2]&A[1]&B[0]&c0)|(B[3]&B[2]&B[1]&A[0]&B[0])|(B[3]&B[2]&B[1]&A[0]&c0)|(B[3]&B[2]&B[1]&B[0]&c0);
assign c5 = (A[4]&B[4])|(A[4]&A[3]&B[3])|(A[4]&A[3]&A[2]&B[2])|(A[4]&A[3]&A[2]&A[1]&B[1])|(A[4]&A[3]&A[2]&A[1]&A[0]&B[0])|(A[4]&A[3]&A[2]&A[1]&A[0]&c0)|(A[4]&A[3]&A[2]&A[1]&B[0]&c0)|(A[4]&A[3]&A[2]&B[1]&A[0]&B[0])|(A[4]&A[3]&A[2]&B[1]&A[0]&c0)|(A[4]&A[3]&A[2]&B[1]&B[0]&c0)|(A[4]&A[3]&B[2]&A[1]&B[1])|(A[4]&A[3]&B[2]&A[1]&A[0]&B[0])|(A[4]&A[3]&B[2]&A[1]&A[0]&c0)|(A[4]&A[3]&B[2]&A[1]&B[0]&c0)|(A[4]&A[3]&B[2]&B[1]&A[0]&B[0])|(A[4]&A[3]&B[2]&B[1]&A[0]&c0)|(A[4]&A[3]&B[2]&B[1]&B[0]&c0)|(A[4]&B[3]&A[2]&B[2])|(A[4]&B[3]&A[2]&A[1]&B[1])|(A[4]&B[3]&A[2]&A[1]&A[0]&B[0])|(A[4]&B[3]&A[2]&A[1]&A[0]&c0)|(A[4]&B[3]&A[2]&A[1]&B[0]&c0)|(A[4]&B[3]&A[2]&B[1]&A[0]&B[0])|(A[4]&B[3]&A[2]&B[1]&A[0]&c0)|(A[4]&B[3]&A[2]&B[1]&B[0]&c0)|(A[4]&B[3]&B[2]&A[1]&B[1])|(A[4]&B[3]&B[2]&A[1]&A[0]&B[0])|(A[4]&B[3]&B[2]&A[1]&A[0]&c0)|(A[4]&B[3]&B[2]&A[1]&B[0]&c0)|(A[4]&B[3]&B[2]&B[1]&A[0]&B[0])|(A[4]&B[3]&B[2]&B[1]&A[0]&c0)|(A[4]&B[3]&B[2]&B[1]&B[0]&c0)|(B[4]&A[3]&B[3])|(B[4]&A[3]&A[2]&B[2])|(B[4]&A[3]&A[2]&A[1]&B[1])|(B[4]&A[3]&A[2]&A[1]&A[0]&B[0])|(B[4]&A[3]&A[2]&A[1]&A[0]&c0)|(B[4]&A[3]&A[2]&A[1]&B[0]&c0)|(B[4]&A[3]&A[2]&B[1]&A[0]&B[0])|(B[4]&A[3]&A[2]&B[1]&A[0]&c0)|(B[4]&A[3]&A[2]&B[1]&B[0]&c0)|(B[4]&A[3]&B[2]&A[1]&B[1])|(B[4]&A[3]&B[2]&A[1]&A[0]&B[0])|(B[4]&A[3]&B[2]&A[1]&A[0]&c0)|(B[4]&A[3]&B[2]&A[1]&B[0]&c0)|(B[4]&A[3]&B[2]&B[1]&A[0]&B[0])|(B[4]&A[3]&B[2]&B[1]&A[0]&c0)|(B[4]&A[3]&B[2]&B[1]&B[0]&c0)|(B[4]&B[3]&A[2]&B[2])|(B[4]&B[3]&A[2]&A[1]&B[1])|(B[4]&B[3]&A[2]&A[1]&A[0]&B[0])|(B[4]&B[3]&A[2]&A[1]&A[0]&c0)|(B[4]&B[3]&A[2]&A[1]&B[0]&c0)|(B[4]&B[3]&A[2]&B[1]&A[0]&B[0])|(B[4]&B[3]&A[2]&B[1]&A[0]&c0)|(B[4]&B[3]&A[2]&B[1]&B[0]&c0)|(B[4]&B[3]&B[2]&A[1]&B[1])|(B[4]&B[3]&B[2]&A[1]&A[0]&B[0])|(B[4]&B[3]&B[2]&A[1]&A[0]&c0)|(B[4]&B[3]&B[2]&A[1]&B[0]&c0)|(B[4]&B[3]&B[2]&B[1]&A[0]&B[0])|(B[4]&B[3]&B[2]&B[1]&A[0]&c0)|(B[4]&B[3]&B[2]&B[1]&B[0]&c0);
assign c6 = (A[5]&B[5])|(A[5]&A[4]&B[4])|(A[5]&A[4]&A[3]&B[3])|(A[5]&A[4]&A[3]&A[2]&B[2])|(A[5]&A[4]&A[3]&A[2]&A[1]&B[1])|(A[5]&A[4]&A[3]&A[2]&A[1]&A[0]&B[0])|(A[5]&A[4]&A[3]&A[2]&A[1]&A[0]&c0)|(A[5]&A[4]&A[3]&A[2]&A[1]&B[0]&c0)|(A[5]&A[4]&A[3]&A[2]&B[1]&A[0]&B[0])|(A[5]&A[4]&A[3]&A[2]&B[1]&A[0]&c0)|(A[5]&A[4]&A[3]&A[2]&B[1]&B[0]&c0)|(A[5]&A[4]&A[3]&B[2]&A[1]&B[1])|(A[5]&A[4]&A[3]&B[2]&A[1]&A[0]&B[0])|(A[5]&A[4]&A[3]&B[2]&A[1]&A[0]&c0)|(A[5]&A[4]&A[3]&B[2]&A[1]&B[0]&c0)|(A[5]&A[4]&A[3]&B[2]&B[1]&A[0]&B[0])|(A[5]&A[4]&A[3]&B[2]&B[1]&A[0]&c0)|(A[5]&A[4]&A[3]&B[2]&B[1]&B[0]&c0)|(A[5]&A[4]&B[3]&A[2]&B[2])|(A[5]&A[4]&B[3]&A[2]&A[1]&B[1])|(A[5]&A[4]&B[3]&A[2]&A[1]&A[0]&B[0])|(A[5]&A[4]&B[3]&A[2]&A[1]&A[0]&c0)|(A[5]&A[4]&B[3]&A[2]&A[1]&B[0]&c0)|(A[5]&A[4]&B[3]&A[2]&B[1]&A[0]&B[0])|(A[5]&A[4]&B[3]&A[2]&B[1]&A[0]&c0)|(A[5]&A[4]&B[3]&A[2]&B[1]&B[0]&c0)|(A[5]&A[4]&B[3]&B[2]&A[1]&B[1])|(A[5]&A[4]&B[3]&B[2]&A[1]&A[0]&B[0])|(A[5]&A[4]&B[3]&B[2]&A[1]&A[0]&c0)|(A[5]&A[4]&B[3]&B[2]&A[1]&B[0]&c0)|(A[5]&A[4]&B[3]&B[2]&B[1]&A[0]&B[0])|(A[5]&A[4]&B[3]&B[2]&B[1]&A[0]&c0)|(A[5]&A[4]&B[3]&B[2]&B[1]&B[0]&c0)|(A[5]&B[4]&A[3]&B[3])|(A[5]&B[4]&A[3]&A[2]&B[2])|(A[5]&B[4]&A[3]&A[2]&A[1]&B[1])|(A[5]&B[4]&A[3]&A[2]&A[1]&A[0]&B[0])|(A[5]&B[4]&A[3]&A[2]&A[1]&A[0]&c0)|(A[5]&B[4]&A[3]&A[2]&A[1]&B[0]&c0)|(A[5]&B[4]&A[3]&A[2]&B[1]&A[0]&B[0])|(A[5]&B[4]&A[3]&A[2]&B[1]&A[0]&c0)|(A[5]&B[4]&A[3]&A[2]&B[1]&B[0]&c0)|(A[5]&B[4]&A[3]&B[2]&A[1]&B[1])|(A[5]&B[4]&A[3]&B[2]&A[1]&A[0]&B[0])|(A[5]&B[4]&A[3]&B[2]&A[1]&A[0]&c0)|(A[5]&B[4]&A[3]&B[2]&A[1]&B[0]&c0)|(A[5]&B[4]&A[3]&B[2]&B[1]&A[0]&B[0])|(A[5]&B[4]&A[3]&B[2]&B[1]&A[0]&c0)|(A[5]&B[4]&A[3]&B[2]&B[1]&B[0]&c0)|(A[5]&B[4]&B[3]&A[2]&B[2])|(A[5]&B[4]&B[3]&A[2]&A[1]&B[1])|(A[5]&B[4]&B[3]&A[2]&A[1]&A[0]&B[0])|(A[5]&B[4]&B[3]&A[2]&A[1]&A[0]&c0)|(A[5]&B[4]&B[3]&A[2]&A[1]&B[0]&c0)|(A[5]&B[4]&B[3]&A[2]&B[1]&A[0]&B[0])|(A[5]&B[4]&B[3]&A[2]&B[1]&A[0]&c0)|(A[5]&B[4]&B[3]&A[2]&B[1]&B[0]&c0)|(A[5]&B[4]&B[3]&B[2]&A[1]&B[1])|(A[5]&B[4]&B[3]&B[2]&A[1]&A[0]&B[0])|(A[5]&B[4]&B[3]&B[2]&A[1]&A[0]&c0)|(A[5]&B[4]&B[3]&B[2]&A[1]&B[0]&c0)|(A[5]&B[4]&B[3]&B[2]&B[1]&A[0]&B[0])|(A[5]&B[4]&B[3]&B[2]&B[1]&A[0]&c0)|(A[5]&B[4]&B[3]&B[2]&B[1]&B[0]&c0)|(B[5]&A[4]&B[4])|(B[5]&A[4]&A[3]&B[3])|(B[5]&A[4]&A[3]&A[2]&B[2])|(B[5]&A[4]&A[3]&A[2]&A[1]&B[1])|(B[5]&A[4]&A[3]&A[2]&A[1]&A[0]&B[0])|(B[5]&A[4]&A[3]&A[2]&A[1]&A[0]&c0)|(B[5]&A[4]&A[3]&A[2]&A[1]&B[0]&c0)|(B[5]&A[4]&A[3]&A[2]&B[1]&A[0]&B[0])|(B[5]&A[4]&A[3]&A[2]&B[1]&A[0]&c0)|(B[5]&A[4]&A[3]&A[2]&B[1]&B[0]&c0)|(B[5]&A[4]&A[3]&B[2]&A[1]&B[1])|(B[5]&A[4]&A[3]&B[2]&A[1]&A[0]&B[0])|(B[5]&A[4]&A[3]&B[2]&A[1]&A[0]&c0)|(B[5]&A[4]&A[3]&B[2]&A[1]&B[0]&c0)|(B[5]&A[4]&A[3]&B[2]&B[1]&A[0]&B[0])|(B[5]&A[4]&A[3]&B[2]&B[1]&A[0]&c0)|(B[5]&A[4]&A[3]&B[2]&B[1]&B[0]&c0)|(B[5]&A[4]&B[3]&A[2]&B[2])|(B[5]&A[4]&B[3]&A[2]&A[1]&B[1])|(B[5]&A[4]&B[3]&A[2]&A[1]&A[0]&B[0])|(B[5]&A[4]&B[3]&A[2]&A[1]&A[0]&c0)|(B[5]&A[4]&B[3]&A[2]&A[1]&B[0]&c0)|(B[5]&A[4]&B[3]&A[2]&B[1]&A[0]&B[0])|(B[5]&A[4]&B[3]&A[2]&B[1]&A[0]&c0)|(B[5]&A[4]&B[3]&A[2]&B[1]&B[0]&c0)|(B[5]&A[4]&B[3]&B[2]&A[1]&B[1])|(B[5]&A[4]&B[3]&B[2]&A[1]&A[0]&B[0])|(B[5]&A[4]&B[3]&B[2]&A[1]&A[0]&c0)|(B[5]&A[4]&B[3]&B[2]&A[1]&B[0]&c0)|(B[5]&A[4]&B[3]&B[2]&B[1]&A[0]&B[0])|(B[5]&A[4]&B[3]&B[2]&B[1]&A[0]&c0)|(B[5]&A[4]&B[3]&B[2]&B[1]&B[0]&c0)|(B[5]&B[4]&A[3]&B[3])|(B[5]&B[4]&A[3]&A[2]&B[2])|(B[5]&B[4]&A[3]&A[2]&A[1]&B[1])|(B[5]&B[4]&A[3]&A[2]&A[1]&A[0]&B[0])|(B[5]&B[4]&A[3]&A[2]&A[1]&A[0]&c0)|(B[5]&B[4]&A[3]&A[2]&A[1]&B[0]&c0)|(B[5]&B[4]&A[3]&A[2]&B[1]&A[0]&B[0])|(B[5]&B[4]&A[3]&A[2]&B[1]&A[0]&c0)|(B[5]&B[4]&A[3]&A[2]&B[1]&B[0]&c0)|(B[5]&B[4]&A[3]&B[2]&A[1]&B[1])|(B[5]&B[4]&A[3]&B[2]&A[1]&A[0]&B[0])|(B[5]&B[4]&A[3]&B[2]&A[1]&A[0]&c0)|(B[5]&B[4]&A[3]&B[2]&A[1]&B[0]&c0)|(B[5]&B[4]&A[3]&B[2]&B[1]&A[0]&B[0])|(B[5]&B[4]&A[3]&B[2]&B[1]&A[0]&c0)|(B[5]&B[4]&A[3]&B[2]&B[1]&B[0]&c0)|(B[5]&B[4]&B[3]&A[2]&B[2])|(B[5]&B[4]&B[3]&A[2]&A[1]&B[1])|(B[5]&B[4]&B[3]&A[2]&A[1]&A[0]&B[0])|(B[5]&B[4]&B[3]&A[2]&A[1]&A[0]&c0)|(B[5]&B[4]&B[3]&A[2]&A[1]&B[0]&c0)|(B[5]&B[4]&B[3]&A[2]&B[1]&A[0]&B[0])|(B[5]&B[4]&B[3]&A[2]&B[1]&A[0]&c0)|(B[5]&B[4]&B[3]&A[2]&B[1]&B[0]&c0)|(B[5]&B[4]&B[3]&B[2]&A[1]&B[1])|(B[5]&B[4]&B[3]&B[2]&A[1]&A[0]&B[0])|(B[5]&B[4]&B[3]&B[2]&A[1]&A[0]&c0)|(B[5]&B[4]&B[3]&B[2]&A[1]&B[0]&c0)|(B[5]&B[4]&B[3]&B[2]&B[1]&A[0]&B[0])|(B[5]&B[4]&B[3]&B[2]&B[1]&A[0]&c0)|(B[5]&B[4]&B[3]&B[2]&B[1]&B[0]&c0);




assign R[0] = A[0] ^ B[0] ^ c0;
assign R[1] = A[1] ^ B[1] ^ c1;
assign R[2] = A[2] ^ B[2] ^ c2;
assign R[3] = A[3] ^ B[3] ^ c3;
assign R[4] = A[4] ^ B[4] ^ c4;
assign R[5] = A[5] ^ B[5] ^ c5;
assign R[6] = A[6] ^ B[6] ^ c6;

endmodule
