module Reg128
(
input [6:0] Rd_Addr, Rs_Addr, Rm_Addr,
input Rd_Wen, Rs_Wen,
input [15:0] Rd_Data, Rs_Data,

output [15:0] Rd_Out, Rs_Out, Rm_Out,

input Clock

);
// the 128 registers
reg [15:0] R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15,R16,R17,R18,R19,R20,R21,R22,R23,R24,R25,R26,R27,R28,R29,R30,R31,R32,R33,R34,R35,R36,R37,R38,R39,R40,R41,R42,R43,R44,R45,R46,R47,R48,R49,R50,R51,R52,R53,R54,R55,R56,R57,R58,R59,R60,R61,R62,R63,R64,R65,R66,R67,R68,R69,R70,R71,R72,R73,R74,R75,R76,R77,R78,R79,R80,R81,R82,R83,R84,R85,R86,R87,R88,R89,R90,R91,R92,R93,R94,R95,R96,R97,R98,R99,R100,R101,R102,R103,R104,R105,R106,R107,R108,R109,R110,R111,R112,R113,R114,R115,R116,R117,R118,R119,R120,R121,R122,R123,R124,R125,R126,R127;
reg [15:0] RdOut, RsOut, RmOut;
assign Rd_Out = RdOut;
assign Rs_Out = RsOut;
assign Rm_Out = RmOut;


// To read data without clock
always @(*) begin
    case(Rd_Addr)
        7'd0 : RdOut = R0;
        7'd1 : RdOut = R1;
        7'd2 : RdOut = R2;
        7'd3 : RdOut = R3;
        7'd4 : RdOut = R4;
        7'd5 : RdOut = R5;
        7'd6 : RdOut = R6;
        7'd7 : RdOut = R7;
        7'd8 : RdOut = R8;
        7'd9 : RdOut = R9;
        7'd10 : RdOut = R10;
        7'd11 : RdOut = R11;
        7'd12 : RdOut = R12;
        7'd13 : RdOut = R13;
        7'd14 : RdOut = R14;
        7'd15 : RdOut = R15;
        7'd16 : RdOut = R16;
        7'd17 : RdOut = R17;
        7'd18 : RdOut = R18;
        7'd19 : RdOut = R19;
        7'd20 : RdOut = R20;
        7'd21 : RdOut = R21;
        7'd22 : RdOut = R22;
        7'd23 : RdOut = R23;
        7'd24 : RdOut = R24;
        7'd25 : RdOut = R25;
        7'd26 : RdOut = R26;
        7'd27 : RdOut = R27;
        7'd28 : RdOut = R28;
        7'd29 : RdOut = R29;
        7'd30 : RdOut = R30;
        7'd31 : RdOut = R31;
        7'd32 : RdOut = R32;
        7'd33 : RdOut = R33;
        7'd34 : RdOut = R34;
        7'd35 : RdOut = R35;
        7'd36 : RdOut = R36;
        7'd37 : RdOut = R37;
        7'd38 : RdOut = R38;
        7'd39 : RdOut = R39;
        7'd40 : RdOut = R40;
        7'd41 : RdOut = R41;
        7'd42 : RdOut = R42;
        7'd43 : RdOut = R43;
        7'd44 : RdOut = R44;
        7'd45 : RdOut = R45;
        7'd46 : RdOut = R46;
        7'd47 : RdOut = R47;
        7'd48 : RdOut = R48;
        7'd49 : RdOut = R49;
        7'd50 : RdOut = R50;
        7'd51 : RdOut = R51;
        7'd52 : RdOut = R52;
        7'd53 : RdOut = R53;
        7'd54 : RdOut = R54;
        7'd55 : RdOut = R55;
        7'd56 : RdOut = R56;
        7'd57 : RdOut = R57;
        7'd58 : RdOut = R58;
        7'd59 : RdOut = R59;
        7'd60 : RdOut = R60;
        7'd61 : RdOut = R61;
        7'd62 : RdOut = R62;
        7'd63 : RdOut = R63;
        7'd64 : RdOut = R64;
        7'd65 : RdOut = R65;
        7'd66 : RdOut = R66;
        7'd67 : RdOut = R67;
        7'd68 : RdOut = R68;
        7'd69 : RdOut = R69;
        7'd70 : RdOut = R70;
        7'd71 : RdOut = R71;
        7'd72 : RdOut = R72;
        7'd73 : RdOut = R73;
        7'd74 : RdOut = R74;
        7'd75 : RdOut = R75;
        7'd76 : RdOut = R76;
        7'd77 : RdOut = R77;
        7'd78 : RdOut = R78;
        7'd79 : RdOut = R79;
        7'd80 : RdOut = R80;
        7'd81 : RdOut = R81;
        7'd82 : RdOut = R82;
        7'd83 : RdOut = R83;
        7'd84 : RdOut = R84;
        7'd85 : RdOut = R85;
        7'd86 : RdOut = R86;
        7'd87 : RdOut = R87;
        7'd88 : RdOut = R88;
        7'd89 : RdOut = R89;
        7'd90 : RdOut = R90;
        7'd91 : RdOut = R91;
        7'd92 : RdOut = R92;
        7'd93 : RdOut = R93;
        7'd94 : RdOut = R94;
        7'd95 : RdOut = R95;
        7'd96 : RdOut = R96;
        7'd97 : RdOut = R97;
        7'd98 : RdOut = R98;
        7'd99 : RdOut = R99;
        7'd100 : RdOut = R100;
        7'd101 : RdOut = R101;
        7'd102 : RdOut = R102;
        7'd103 : RdOut = R103;
        7'd104 : RdOut = R104;
        7'd105 : RdOut = R105;
        7'd106 : RdOut = R106;
        7'd107 : RdOut = R107;
        7'd108 : RdOut = R108;
        7'd109 : RdOut = R109;
        7'd110 : RdOut = R110;
        7'd111 : RdOut = R111;
        7'd112 : RdOut = R112;
        7'd113 : RdOut = R113;
        7'd114 : RdOut = R114;
        7'd115 : RdOut = R115;
        7'd116 : RdOut = R116;
        7'd117 : RdOut = R117;
        7'd118 : RdOut = R118;
        7'd119 : RdOut = R119;
        7'd120 : RdOut = R120;
        7'd121 : RdOut = R121;
        7'd122 : RdOut = R122;
        7'd123 : RdOut = R123;
        7'd124 : RdOut = R124;
        7'd125 : RdOut = R125;
        7'd126 : RdOut = R126;
        7'd127 : RdOut = R127;

    endcase

    case(Rs_Addr)
        7'd0 : RsOut = R0;
        7'd1 : RsOut = R1;
        7'd2 : RsOut = R2;
        7'd3 : RsOut = R3;
        7'd4 : RsOut = R4;
        7'd5 : RsOut = R5;
        7'd6 : RsOut = R6;
        7'd7 : RsOut = R7;
        7'd8 : RsOut = R8;
        7'd9 : RsOut = R9;
        7'd10 : RsOut = R10;
        7'd11 : RsOut = R11;
        7'd12 : RsOut = R12;
        7'd13 : RsOut = R13;
        7'd14 : RsOut = R14;
        7'd15 : RsOut = R15;
        7'd16 : RsOut = R16;
        7'd17 : RsOut = R17;
        7'd18 : RsOut = R18;
        7'd19 : RsOut = R19;
        7'd20 : RsOut = R20;
        7'd21 : RsOut = R21;
        7'd22 : RsOut = R22;
        7'd23 : RsOut = R23;
        7'd24 : RsOut = R24;
        7'd25 : RsOut = R25;
        7'd26 : RsOut = R26;
        7'd27 : RsOut = R27;
        7'd28 : RsOut = R28;
        7'd29 : RsOut = R29;
        7'd30 : RsOut = R30;
        7'd31 : RsOut = R31;
        7'd32 : RsOut = R32;
        7'd33 : RsOut = R33;
        7'd34 : RsOut = R34;
        7'd35 : RsOut = R35;
        7'd36 : RsOut = R36;
        7'd37 : RsOut = R37;
        7'd38 : RsOut = R38;
        7'd39 : RsOut = R39;
        7'd40 : RsOut = R40;
        7'd41 : RsOut = R41;
        7'd42 : RsOut = R42;
        7'd43 : RsOut = R43;
        7'd44 : RsOut = R44;
        7'd45 : RsOut = R45;
        7'd46 : RsOut = R46;
        7'd47 : RsOut = R47;
        7'd48 : RsOut = R48;
        7'd49 : RsOut = R49;
        7'd50 : RsOut = R50;
        7'd51 : RsOut = R51;
        7'd52 : RsOut = R52;
        7'd53 : RsOut = R53;
        7'd54 : RsOut = R54;
        7'd55 : RsOut = R55;
        7'd56 : RsOut = R56;
        7'd57 : RsOut = R57;
        7'd58 : RsOut = R58;
        7'd59 : RsOut = R59;
        7'd60 : RsOut = R60;
        7'd61 : RsOut = R61;
        7'd62 : RsOut = R62;
        7'd63 : RsOut = R63;
        7'd64 : RsOut = R64;
        7'd65 : RsOut = R65;
        7'd66 : RsOut = R66;
        7'd67 : RsOut = R67;
        7'd68 : RsOut = R68;
        7'd69 : RsOut = R69;
        7'd70 : RsOut = R70;
        7'd71 : RsOut = R71;
        7'd72 : RsOut = R72;
        7'd73 : RsOut = R73;
        7'd74 : RsOut = R74;
        7'd75 : RsOut = R75;
        7'd76 : RsOut = R76;
        7'd77 : RsOut = R77;
        7'd78 : RsOut = R78;
        7'd79 : RsOut = R79;
        7'd80 : RsOut = R80;
        7'd81 : RsOut = R81;
        7'd82 : RsOut = R82;
        7'd83 : RsOut = R83;
        7'd84 : RsOut = R84;
        7'd85 : RsOut = R85;
        7'd86 : RsOut = R86;
        7'd87 : RsOut = R87;
        7'd88 : RsOut = R88;
        7'd89 : RsOut = R89;
        7'd90 : RsOut = R90;
        7'd91 : RsOut = R91;
        7'd92 : RsOut = R92;
        7'd93 : RsOut = R93;
        7'd94 : RsOut = R94;
        7'd95 : RsOut = R95;
        7'd96 : RsOut = R96;
        7'd97 : RsOut = R97;
        7'd98 : RsOut = R98;
        7'd99 : RsOut = R99;
        7'd100 : RsOut = R100;
        7'd101 : RsOut = R101;
        7'd102 : RsOut = R102;
        7'd103 : RsOut = R103;
        7'd104 : RsOut = R104;
        7'd105 : RsOut = R105;
        7'd106 : RsOut = R106;
        7'd107 : RsOut = R107;
        7'd108 : RsOut = R108;
        7'd109 : RsOut = R109;
        7'd110 : RsOut = R110;
        7'd111 : RsOut = R111;
        7'd112 : RsOut = R112;
        7'd113 : RsOut = R113;
        7'd114 : RsOut = R114;
        7'd115 : RsOut = R115;
        7'd116 : RsOut = R116;
        7'd117 : RsOut = R117;
        7'd118 : RsOut = R118;
        7'd119 : RsOut = R119;
        7'd120 : RsOut = R120;
        7'd121 : RsOut = R121;
        7'd122 : RsOut = R122;
        7'd123 : RsOut = R123;
        7'd124 : RsOut = R124;
        7'd125 : RsOut = R125;
        7'd126 : RsOut = R126;
        7'd127 : RsOut = R127;

    endcase

    case(Rm_Addr)
        7'd0 : RmOut = R0;
        7'd1 : RmOut = R1;
        7'd2 : RmOut = R2;
        7'd3 : RmOut = R3;
        7'd4 : RmOut = R4;
        7'd5 : RmOut = R5;
        7'd6 : RmOut = R6;
        7'd7 : RmOut = R7;
        7'd8 : RmOut = R8;
        7'd9 : RmOut = R9;
        7'd10 : RmOut = R10;
        7'd11 : RmOut = R11;
        7'd12 : RmOut = R12;
        7'd13 : RmOut = R13;
        7'd14 : RmOut = R14;
        7'd15 : RmOut = R15;
        7'd16 : RmOut = R16;
        7'd17 : RmOut = R17;
        7'd18 : RmOut = R18;
        7'd19 : RmOut = R19;
        7'd20 : RmOut = R20;
        7'd21 : RmOut = R21;
        7'd22 : RmOut = R22;
        7'd23 : RmOut = R23;
        7'd24 : RmOut = R24;
        7'd25 : RmOut = R25;
        7'd26 : RmOut = R26;
        7'd27 : RmOut = R27;
        7'd28 : RmOut = R28;
        7'd29 : RmOut = R29;
        7'd30 : RmOut = R30;
        7'd31 : RmOut = R31;
        7'd32 : RmOut = R32;
        7'd33 : RmOut = R33;
        7'd34 : RmOut = R34;
        7'd35 : RmOut = R35;
        7'd36 : RmOut = R36;
        7'd37 : RmOut = R37;
        7'd38 : RmOut = R38;
        7'd39 : RmOut = R39;
        7'd40 : RmOut = R40;
        7'd41 : RmOut = R41;
        7'd42 : RmOut = R42;
        7'd43 : RmOut = R43;
        7'd44 : RmOut = R44;
        7'd45 : RmOut = R45;
        7'd46 : RmOut = R46;
        7'd47 : RmOut = R47;
        7'd48 : RmOut = R48;
        7'd49 : RmOut = R49;
        7'd50 : RmOut = R50;
        7'd51 : RmOut = R51;
        7'd52 : RmOut = R52;
        7'd53 : RmOut = R53;
        7'd54 : RmOut = R54;
        7'd55 : RmOut = R55;
        7'd56 : RmOut = R56;
        7'd57 : RmOut = R57;
        7'd58 : RmOut = R58;
        7'd59 : RmOut = R59;
        7'd60 : RmOut = R60;
        7'd61 : RmOut = R61;
        7'd62 : RmOut = R62;
        7'd63 : RmOut = R63;
        7'd64 : RmOut = R64;
        7'd65 : RmOut = R65;
        7'd66 : RmOut = R66;
        7'd67 : RmOut = R67;
        7'd68 : RmOut = R68;
        7'd69 : RmOut = R69;
        7'd70 : RmOut = R70;
        7'd71 : RmOut = R71;
        7'd72 : RmOut = R72;
        7'd73 : RmOut = R73;
        7'd74 : RmOut = R74;
        7'd75 : RmOut = R75;
        7'd76 : RmOut = R76;
        7'd77 : RmOut = R77;
        7'd78 : RmOut = R78;
        7'd79 : RmOut = R79;
        7'd80 : RmOut = R80;
        7'd81 : RmOut = R81;
        7'd82 : RmOut = R82;
        7'd83 : RmOut = R83;
        7'd84 : RmOut = R84;
        7'd85 : RmOut = R85;
        7'd86 : RmOut = R86;
        7'd87 : RmOut = R87;
        7'd88 : RmOut = R88;
        7'd89 : RmOut = R89;
        7'd90 : RmOut = R90;
        7'd91 : RmOut = R91;
        7'd92 : RmOut = R92;
        7'd93 : RmOut = R93;
        7'd94 : RmOut = R94;
        7'd95 : RmOut = R95;
        7'd96 : RmOut = R96;
        7'd97 : RmOut = R97;
        7'd98 : RmOut = R98;
        7'd99 : RmOut = R99;
        7'd100 : RmOut = R100;
        7'd101 : RmOut = R101;
        7'd102 : RmOut = R102;
        7'd103 : RmOut = R103;
        7'd104 : RmOut = R104;
        7'd105 : RmOut = R105;
        7'd106 : RmOut = R106;
        7'd107 : RmOut = R107;
        7'd108 : RmOut = R108;
        7'd109 : RmOut = R109;
        7'd110 : RmOut = R110;
        7'd111 : RmOut = R111;
        7'd112 : RmOut = R112;
        7'd113 : RmOut = R113;
        7'd114 : RmOut = R114;
        7'd115 : RmOut = R115;
        7'd116 : RmOut = R116;
        7'd117 : RmOut = R117;
        7'd118 : RmOut = R118;
        7'd119 : RmOut = R119;
        7'd120 : RmOut = R120;
        7'd121 : RmOut = R121;
        7'd122 : RmOut = R122;
        7'd123 : RmOut = R123;
        7'd124 : RmOut = R124;
        7'd125 : RmOut = R125;
        7'd126 : RmOut = R126;
        7'd127 : RmOut = R127;

    endcase
end

// To write data on positive edge of clock
always @(posedge Clock) begin
    if(Rd_Wen)
        case(Rd_Addr)
            7'd0 : R0 <= Rd_Data;
            7'd1 : R1 <= Rd_Data;
            7'd2 : R2 <= Rd_Data;
            7'd3 : R3 <= Rd_Data;
            7'd4 : R4 <= Rd_Data;
            7'd5 : R5 <= Rd_Data;
            7'd6 : R6 <= Rd_Data;
            7'd7 : R7 <= Rd_Data;
            7'd8 : R8 <= Rd_Data;
            7'd9 : R9 <= Rd_Data;
            7'd10 : R10 <= Rd_Data;
            7'd11 : R11 <= Rd_Data;
            7'd12 : R12 <= Rd_Data;
            7'd13 : R13 <= Rd_Data;
            7'd14 : R14 <= Rd_Data;
            7'd15 : R15 <= Rd_Data;
            7'd16 : R16 <= Rd_Data;
            7'd17 : R17 <= Rd_Data;
            7'd18 : R18 <= Rd_Data;
            7'd19 : R19 <= Rd_Data;
            7'd20 : R20 <= Rd_Data;
            7'd21 : R21 <= Rd_Data;
            7'd22 : R22 <= Rd_Data;
            7'd23 : R23 <= Rd_Data;
            7'd24 : R24 <= Rd_Data;
            7'd25 : R25 <= Rd_Data;
            7'd26 : R26 <= Rd_Data;
            7'd27 : R27 <= Rd_Data;
            7'd28 : R28 <= Rd_Data;
            7'd29 : R29 <= Rd_Data;
            7'd30 : R30 <= Rd_Data;
            7'd31 : R31 <= Rd_Data;
            7'd32 : R32 <= Rd_Data;
            7'd33 : R33 <= Rd_Data;
            7'd34 : R34 <= Rd_Data;
            7'd35 : R35 <= Rd_Data;
            7'd36 : R36 <= Rd_Data;
            7'd37 : R37 <= Rd_Data;
            7'd38 : R38 <= Rd_Data;
            7'd39 : R39 <= Rd_Data;
            7'd40 : R40 <= Rd_Data;
            7'd41 : R41 <= Rd_Data;
            7'd42 : R42 <= Rd_Data;
            7'd43 : R43 <= Rd_Data;
            7'd44 : R44 <= Rd_Data;
            7'd45 : R45 <= Rd_Data;
            7'd46 : R46 <= Rd_Data;
            7'd47 : R47 <= Rd_Data;
            7'd48 : R48 <= Rd_Data;
            7'd49 : R49 <= Rd_Data;
            7'd50 : R50 <= Rd_Data;
            7'd51 : R51 <= Rd_Data;
            7'd52 : R52 <= Rd_Data;
            7'd53 : R53 <= Rd_Data;
            7'd54 : R54 <= Rd_Data;
            7'd55 : R55 <= Rd_Data;
            7'd56 : R56 <= Rd_Data;
            7'd57 : R57 <= Rd_Data;
            7'd58 : R58 <= Rd_Data;
            7'd59 : R59 <= Rd_Data;
            7'd60 : R60 <= Rd_Data;
            7'd61 : R61 <= Rd_Data;
            7'd62 : R62 <= Rd_Data;
            7'd63 : R63 <= Rd_Data;
            7'd64 : R64 <= Rd_Data;
            7'd65 : R65 <= Rd_Data;
            7'd66 : R66 <= Rd_Data;
            7'd67 : R67 <= Rd_Data;
            7'd68 : R68 <= Rd_Data;
            7'd69 : R69 <= Rd_Data;
            7'd70 : R70 <= Rd_Data;
            7'd71 : R71 <= Rd_Data;
            7'd72 : R72 <= Rd_Data;
            7'd73 : R73 <= Rd_Data;
            7'd74 : R74 <= Rd_Data;
            7'd75 : R75 <= Rd_Data;
            7'd76 : R76 <= Rd_Data;
            7'd77 : R77 <= Rd_Data;
            7'd78 : R78 <= Rd_Data;
            7'd79 : R79 <= Rd_Data;
            7'd80 : R80 <= Rd_Data;
            7'd81 : R81 <= Rd_Data;
            7'd82 : R82 <= Rd_Data;
            7'd83 : R83 <= Rd_Data;
            7'd84 : R84 <= Rd_Data;
            7'd85 : R85 <= Rd_Data;
            7'd86 : R86 <= Rd_Data;
            7'd87 : R87 <= Rd_Data;
            7'd88 : R88 <= Rd_Data;
            7'd89 : R89 <= Rd_Data;
            7'd90 : R90 <= Rd_Data;
            7'd91 : R91 <= Rd_Data;
            7'd92 : R92 <= Rd_Data;
            7'd93 : R93 <= Rd_Data;
            7'd94 : R94 <= Rd_Data;
            7'd95 : R95 <= Rd_Data;
            7'd96 : R96 <= Rd_Data;
            7'd97 : R97 <= Rd_Data;
            7'd98 : R98 <= Rd_Data;
            7'd99 : R99 <= Rd_Data;
            7'd100 : R100 <= Rd_Data;
            7'd101 : R101 <= Rd_Data;
            7'd102 : R102 <= Rd_Data;
            7'd103 : R103 <= Rd_Data;
            7'd104 : R104 <= Rd_Data;
            7'd105 : R105 <= Rd_Data;
            7'd106 : R106 <= Rd_Data;
            7'd107 : R107 <= Rd_Data;
            7'd108 : R108 <= Rd_Data;
            7'd109 : R109 <= Rd_Data;
            7'd110 : R110 <= Rd_Data;
            7'd111 : R111 <= Rd_Data;
            7'd112 : R112 <= Rd_Data;
            7'd113 : R113 <= Rd_Data;
            7'd114 : R114 <= Rd_Data;
            7'd115 : R115 <= Rd_Data;
            7'd116 : R116 <= Rd_Data;
            7'd117 : R117 <= Rd_Data;
            7'd118 : R118 <= Rd_Data;
            7'd119 : R119 <= Rd_Data;
            7'd120 : R120 <= Rd_Data;
            7'd121 : R121 <= Rd_Data;
            7'd122 : R122 <= Rd_Data;
            7'd123 : R123 <= Rd_Data;
            7'd124 : R124 <= Rd_Data;
            7'd125 : R125 <= Rd_Data;
            7'd126 : R126 <= Rd_Data;
            7'd127 : R127 <= Rd_Data;
        endcase
    
    if(Rs_Wen)
        case(Rs_Addr)
            7'd0 : R0 <= Rs_Data;
            7'd1 : R1 <= Rs_Data;
            7'd2 : R2 <= Rs_Data;
            7'd3 : R3 <= Rs_Data;
            7'd4 : R4 <= Rs_Data;
            7'd5 : R5 <= Rs_Data;
            7'd6 : R6 <= Rs_Data;
            7'd7 : R7 <= Rs_Data;
            7'd8 : R8 <= Rs_Data;
            7'd9 : R9 <= Rs_Data;
            7'd10 : R10 <= Rs_Data;
            7'd11 : R11 <= Rs_Data;
            7'd12 : R12 <= Rs_Data;
            7'd13 : R13 <= Rs_Data;
            7'd14 : R14 <= Rs_Data;
            7'd15 : R15 <= Rs_Data;
            7'd16 : R16 <= Rs_Data;
            7'd17 : R17 <= Rs_Data;
            7'd18 : R18 <= Rs_Data;
            7'd19 : R19 <= Rs_Data;
            7'd20 : R20 <= Rs_Data;
            7'd21 : R21 <= Rs_Data;
            7'd22 : R22 <= Rs_Data;
            7'd23 : R23 <= Rs_Data;
            7'd24 : R24 <= Rs_Data;
            7'd25 : R25 <= Rs_Data;
            7'd26 : R26 <= Rs_Data;
            7'd27 : R27 <= Rs_Data;
            7'd28 : R28 <= Rs_Data;
            7'd29 : R29 <= Rs_Data;
            7'd30 : R30 <= Rs_Data;
            7'd31 : R31 <= Rs_Data;
            7'd32 : R32 <= Rs_Data;
            7'd33 : R33 <= Rs_Data;
            7'd34 : R34 <= Rs_Data;
            7'd35 : R35 <= Rs_Data;
            7'd36 : R36 <= Rs_Data;
            7'd37 : R37 <= Rs_Data;
            7'd38 : R38 <= Rs_Data;
            7'd39 : R39 <= Rs_Data;
            7'd40 : R40 <= Rs_Data;
            7'd41 : R41 <= Rs_Data;
            7'd42 : R42 <= Rs_Data;
            7'd43 : R43 <= Rs_Data;
            7'd44 : R44 <= Rs_Data;
            7'd45 : R45 <= Rs_Data;
            7'd46 : R46 <= Rs_Data;
            7'd47 : R47 <= Rs_Data;
            7'd48 : R48 <= Rs_Data;
            7'd49 : R49 <= Rs_Data;
            7'd50 : R50 <= Rs_Data;
            7'd51 : R51 <= Rs_Data;
            7'd52 : R52 <= Rs_Data;
            7'd53 : R53 <= Rs_Data;
            7'd54 : R54 <= Rs_Data;
            7'd55 : R55 <= Rs_Data;
            7'd56 : R56 <= Rs_Data;
            7'd57 : R57 <= Rs_Data;
            7'd58 : R58 <= Rs_Data;
            7'd59 : R59 <= Rs_Data;
            7'd60 : R60 <= Rs_Data;
            7'd61 : R61 <= Rs_Data;
            7'd62 : R62 <= Rs_Data;
            7'd63 : R63 <= Rs_Data;
            7'd64 : R64 <= Rs_Data;
            7'd65 : R65 <= Rs_Data;
            7'd66 : R66 <= Rs_Data;
            7'd67 : R67 <= Rs_Data;
            7'd68 : R68 <= Rs_Data;
            7'd69 : R69 <= Rs_Data;
            7'd70 : R70 <= Rs_Data;
            7'd71 : R71 <= Rs_Data;
            7'd72 : R72 <= Rs_Data;
            7'd73 : R73 <= Rs_Data;
            7'd74 : R74 <= Rs_Data;
            7'd75 : R75 <= Rs_Data;
            7'd76 : R76 <= Rs_Data;
            7'd77 : R77 <= Rs_Data;
            7'd78 : R78 <= Rs_Data;
            7'd79 : R79 <= Rs_Data;
            7'd80 : R80 <= Rs_Data;
            7'd81 : R81 <= Rs_Data;
            7'd82 : R82 <= Rs_Data;
            7'd83 : R83 <= Rs_Data;
            7'd84 : R84 <= Rs_Data;
            7'd85 : R85 <= Rs_Data;
            7'd86 : R86 <= Rs_Data;
            7'd87 : R87 <= Rs_Data;
            7'd88 : R88 <= Rs_Data;
            7'd89 : R89 <= Rs_Data;
            7'd90 : R90 <= Rs_Data;
            7'd91 : R91 <= Rs_Data;
            7'd92 : R92 <= Rs_Data;
            7'd93 : R93 <= Rs_Data;
            7'd94 : R94 <= Rs_Data;
            7'd95 : R95 <= Rs_Data;
            7'd96 : R96 <= Rs_Data;
            7'd97 : R97 <= Rs_Data;
            7'd98 : R98 <= Rs_Data;
            7'd99 : R99 <= Rs_Data;
            7'd100 : R100 <= Rs_Data;
            7'd101 : R101 <= Rs_Data;
            7'd102 : R102 <= Rs_Data;
            7'd103 : R103 <= Rs_Data;
            7'd104 : R104 <= Rs_Data;
            7'd105 : R105 <= Rs_Data;
            7'd106 : R106 <= Rs_Data;
            7'd107 : R107 <= Rs_Data;
            7'd108 : R108 <= Rs_Data;
            7'd109 : R109 <= Rs_Data;
            7'd110 : R110 <= Rs_Data;
            7'd111 : R111 <= Rs_Data;
            7'd112 : R112 <= Rs_Data;
            7'd113 : R113 <= Rs_Data;
            7'd114 : R114 <= Rs_Data;
            7'd115 : R115 <= Rs_Data;
            7'd116 : R116 <= Rs_Data;
            7'd117 : R117 <= Rs_Data;
            7'd118 : R118 <= Rs_Data;
            7'd119 : R119 <= Rs_Data;
            7'd120 : R120 <= Rs_Data;
            7'd121 : R121 <= Rs_Data;
            7'd122 : R122 <= Rs_Data;
            7'd123 : R123 <= Rs_Data;
            7'd124 : R124 <= Rs_Data;
            7'd125 : R125 <= Rs_Data;
            7'd126 : R126 <= Rs_Data;
            7'd127 : R127 <= Rs_Data;
        endcase
    
end

endmodule