module add1
(
	input [15:0] i,
	output [15:0] o
);

assign o = i + 1'd1;

endmodule